-- MULTIPLEXOR: m <= (NOT (s) AND x) OR (s AND y);
-- s=0, m=x
