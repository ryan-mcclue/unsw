-- archive 3,4,5
-- .jpeg 4 and 5

-- user manual for pin assignments  
-- reference manual also

-- can target entire vectors

-- segment display 1 indicates particular segment is on

-- mcclue-5346008-lab01-part1.qad

-- testbenches is umbrella term for waveform functional/timing simulation etc.
